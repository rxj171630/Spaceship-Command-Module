module testbench;
initial begin
  forever begin
  $display("Hello World");
  $finish;
  end
end
endmodule
